library verilog;
use verilog.vl_types.all;
entity rpn_vlg_vec_tst is
end rpn_vlg_vec_tst;
